module f_not(x,f);
input x;
output f;
assign f = ~x;
endmodule
